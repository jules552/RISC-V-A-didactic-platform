parameter ALU_ADD = 'b0000;
parameter ALU_SUB = 'b0001;
parameter ALU_XOR = 'b0010;
parameter ALU_OR = 'b0011;
parameter ALU_AND = 'b0100;
parameter ALU_SSL = 'b0101;
parameter ALU_SRL = 'b0110;
parameter ALU_SRA = 'b0111;
parameter ALU_SLT = 'b1000;
parameter ALU_SLTU = 'b1001;
parameter ALU_NOP = 'b1010;
parameter ALU_INVALID = 'b1111;